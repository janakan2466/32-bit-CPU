library verilog;
use verilog.vl_types.all;
entity register32_vlg_vec_tst is
end register32_vlg_vec_tst;
