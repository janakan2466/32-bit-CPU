library verilog;
use verilog.vl_types.all;
entity adder32_vlg_vec_tst is
end adder32_vlg_vec_tst;
