library verilog;
use verilog.vl_types.all;
entity mux2to1_vlg_vec_tst is
end mux2to1_vlg_vec_tst;
