library verilog;
use verilog.vl_types.all;
entity CPU_TEST_Sim_vlg_vec_tst is
end CPU_TEST_Sim_vlg_vec_tst;
