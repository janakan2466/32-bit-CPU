library verilog;
use verilog.vl_types.all;
entity Control_New_vlg_vec_tst is
end Control_New_vlg_vec_tst;
