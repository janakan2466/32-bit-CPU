library verilog;
use verilog.vl_types.all;
entity adder4_vlg_vec_tst is
end adder4_vlg_vec_tst;
