library verilog;
use verilog.vl_types.all;
entity data_mem_vlg_vec_tst is
end data_mem_vlg_vec_tst;
