library verilog;
use verilog.vl_types.all;
entity add_vlg_vec_tst is
end add_vlg_vec_tst;
