library verilog;
use verilog.vl_types.all;
entity register1_vlg_vec_tst is
end register1_vlg_vec_tst;
