library verilog;
use verilog.vl_types.all;
entity fulladd_vlg_vec_tst is
end fulladd_vlg_vec_tst;
