library verilog;
use verilog.vl_types.all;
entity ControlUnit_vlg_vec_tst is
end ControlUnit_vlg_vec_tst;
