library verilog;
use verilog.vl_types.all;
entity adder16_vlg_vec_tst is
end adder16_vlg_vec_tst;
