library verilog;
use verilog.vl_types.all;
entity ControlUnit2_vlg_vec_tst is
end ControlUnit2_vlg_vec_tst;
