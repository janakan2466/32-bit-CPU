library verilog;
use verilog.vl_types.all;
entity reset_circuit_vlg_vec_tst is
end reset_circuit_vlg_vec_tst;
