library verilog;
use verilog.vl_types.all;
entity data_path_vlg_vec_tst is
end data_path_vlg_vec_tst;
